// 시스템 컨트롤러 정의
module sc;

endmodule