// 1bit 전가산기(FA)모듈 생성
module fa;

endmodule