// 공유 메모리 모듈 정의
module mem;

endmodule