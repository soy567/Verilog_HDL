// 데이터 Crossbar 정의
module xbar;

endmodule