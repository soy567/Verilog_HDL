`include "IS.v"

module stimulus;
    is is1();
endmodule